2025(S)-AI-138
